`timescale 1ns / 1ps

module VLSU(

    );
    
    
    
endmodule